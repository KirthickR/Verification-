interface intf;
  logic clk;
  logic we;
  logic re;
  logic [3:0]data_in;
  logic [1:0]addr;
  logic [3:0]data_out;
endinterface
  
